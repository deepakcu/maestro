// ethernet_port_interface_0.v

// Generated using ACDS version 12.0 178 at 2012.08.08.17:01:19

`timescale 1 ps / 1 ps
module ethernet_port_interface_0 (
		input  wire        clk,                      //                   clock.clk
		input  wire        reset,                    //                   reset.reset
		input  wire [26:0] control_port_address,     //            control_port.address
		input  wire        control_port_read,        //                        .read
		output wire [31:0] control_port_readdata,    //                        .readdata
		input  wire        control_port_write,       //                        .write
		input  wire [31:0] control_port_writedata,   //                        .writedata
		output wire        control_port_waitrequest, //                        .waitrequest
		input  wire [7:0]  sink_data0,               //   avalon_streaming_sink.data
		output wire        sink_ready0,              //                        .ready
		input  wire        sink_valid0,              //                        .valid
		input  wire [5:0]  sink_error0,              //                        .error
		input  wire        sink_startofpacket0,      //                        .startofpacket
		input  wire        sink_endofpacket0,        //                        .endofpacket
		output wire [7:0]  source_data0,             // avalon_streaming_source.data
		input  wire        source_ready0,            //                        .ready
		output wire        source_valid0,            //                        .valid
		output wire        source_error0,            //                        .error
		output wire        source_startofpacket0,    //                        .startofpacket
		output wire        source_endofpacket0       //                        .endofpacket
	);

	ethernet_port_interface ethernet_port_interface_0_inst (
		.clk                      (clk),                      //                   clock.clk
		.reset                    (reset),                    //                   reset.reset
		.control_port_address     (control_port_address),     //            control_port.address
		.control_port_read        (control_port_read),        //                        .read
		.control_port_readdata    (control_port_readdata),    //                        .readdata
		.control_port_write       (control_port_write),       //                        .write
		.control_port_writedata   (control_port_writedata),   //                        .writedata
		.control_port_waitrequest (control_port_waitrequest), //                        .waitrequest
		.sink_data0               (sink_data0),               //   avalon_streaming_sink.data
		.sink_ready0              (sink_ready0),              //                        .ready
		.sink_valid0              (sink_valid0),              //                        .valid
		.sink_error0              (sink_error0),              //                        .error
		.sink_startofpacket0      (sink_startofpacket0),      //                        .startofpacket
		.sink_endofpacket0        (sink_endofpacket0),        //                        .endofpacket
		.source_data0             (source_data0),             // avalon_streaming_source.data
		.source_ready0            (source_ready0),            //                        .ready
		.source_valid0            (source_valid0),            //                        .valid
		.source_error0            (source_error0),            //                        .error
		.source_startofpacket0    (source_startofpacket0),    //                        .startofpacket
		.source_endofpacket0      (source_endofpacket0)       //                        .endofpacket
	);

endmodule
